** sch_path: /home/alexa/TemporalChip/xschem/projects/Vernier8Bit.sch
**.subckt Vernier8Bit VDD GND IN1 IN2 t0 t7 t1 t2 t3 t4 t5 t6
*.ipin VDD
*.ipin GND
*.ipin IN1
*.ipin IN2
*.opin t0
*.opin t7
*.opin t1
*.opin t2
*.opin t3
*.opin t4
*.opin t5
*.opin t6
x16 t0 IN1 net1 IN2 VDD GND VernierSymbol
x1 t1 t0 net2 net1 VDD GND VernierSymbol
x2 t2 t1 net3 net2 VDD GND VernierSymbol
x3 t3 t2 net7 net3 VDD GND VernierSymbol
x4 t4 t3 net4 net7 VDD GND VernierSymbol
x7 t5 t4 net5 net4 VDD GND VernierSymbol
x8 t6 t5 net6 net5 VDD GND VernierSymbol
x9 t7 t6 net8 net6 VDD GND VernierSymbol
* noconn #net8
**.ends

* expanding   symbol:  VernierSymbol.sym # of pins=6
** sym_path: /home/alexa/TemporalChip/xschem/projects/VernierSymbol.sym
** sch_path: /home/alexa/TemporalChip/xschem/projects/VernierSymbol.sch
.subckt VernierSymbol OUT1 IN1 OUT2 IN2 VDD GND
*.ipin VDD
*.ipin GND
*.ipin IN1
*.ipin IN2
*.opin OUT1
*.opin OUT2
x2 net8 OUT2 0 0 VDD VDD OUT1 sky130_fd_sc_hd__dlxtp_1
x10 net5 GND GND VDD VDD net7 sky130_fd_sc_hd__buf_1
x11 net4 GND GND VDD VDD net5 sky130_fd_sc_hd__buf_1
x12 IN2 GND GND VDD VDD net4 sky130_fd_sc_hd__buf_1
x6 net3 GND GND VDD VDD net6 sky130_fd_sc_hd__buf_1
x7 net2 GND GND VDD VDD net3 sky130_fd_sc_hd__buf_1
x8 net1 GND GND VDD VDD net2 sky130_fd_sc_hd__buf_1
x9 IN1 GND GND VDD VDD net1 sky130_fd_sc_hd__buf_1
x5 net6 GND GND VDD VDD net8 sky130_fd_sc_hd__buf_1
x13 net7 GND GND VDD VDD OUT2 sky130_fd_sc_hd__buf_1
.ends

.GLOBAL GND
.end
