** sch_path: /home/alexa/TemporalChip/xschem/projects/SingleVernier.sch
**.subckt SingleVernier
V1 VIN1 GND PULSE(0 1.8 0n 100p 100p 5n 10n)
V2 VIN2 GND PULSE(0 1.8 0n 100p 100p 5n 10n)
V3 VDD GND 1.8
x2 net12 net11 0 0 VDD VDD VOUT sky130_fd_sc_hd__dlxtp_1
x10 net5 GND GND VDD VDD net10 sky130_fd_sc_hd__buf_1
x11 net4 GND GND VDD VDD net5 sky130_fd_sc_hd__buf_1
x12 VIN2 GND GND VDD VDD net4 sky130_fd_sc_hd__buf_1
x6 net3 GND GND VDD VDD net9 sky130_fd_sc_hd__buf_1
x7 net2 GND GND VDD VDD net3 sky130_fd_sc_hd__buf_1
x8 net1 GND GND VDD VDD net2 sky130_fd_sc_hd__buf_1
x9 VIN1 GND GND VDD VDD net1 sky130_fd_sc_hd__buf_1
x1 net8 GND GND VDD VDD net12 sky130_fd_sc_hd__buf_1
x3 net7 GND GND VDD VDD net8 sky130_fd_sc_hd__buf_1
x4 net6 GND GND VDD VDD net7 sky130_fd_sc_hd__buf_1
x5 net9 GND GND VDD VDD net6 sky130_fd_sc_hd__buf_1
x13 net10 GND GND VDD VDD net11 sky130_fd_sc_hd__buf_1
**** begin user architecture code


.include /home/alexa/open_pdks/sky130/sky130B/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.control
tran 10p 30n
write /home/alexa/chip_design/xschem/simulations/VernierDelay.raw
plot v(VIN1) v(VOUT)
.endc

.options acct list


.lib /usr/local/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends
.GLOBAL GND
.end
