** sch_path: /home/alexa/TemporalChip/xschem/projects/untitled.sch
**.subckt untitled
V1 VIN1 GND PULSE(0 1.8 0n 100p 100p 5n 10n)
V2 VIN2 GND PULSE(0 1.8 0n 100p 100p 5n 10n)
V3 VDD GND 1.8
x2 VIN1 VIN2 0 0 VDD VDD VOUT sky130_fd_sc_hd__dlxtp_1
**** begin user architecture code


.include /home/alexa/open_pdks/sky130/sky130B/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.control
tran 10p 30n
write /home/alexa/chip_design/xschem/simulations/VernierDelay.raw
plot v(VIN1) v(VOUT)
.endc

.options acct list


.lib /usr/local/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends
.GLOBAL GND
.end
