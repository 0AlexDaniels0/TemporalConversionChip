** sch_path: /home/alexa/TemporalChip/xschem/projects/VernierArray.sch
**.subckt VernierArray
V1 VIN2 GND PULSE(0 1.8 0n 100p 100p 5n 20n)
V2 VIN1 GND PULSE(0 1.8 0n 100p 100p 5n 10n)
V3 VDD GND 1.8
x16 net2 VIN1 net1 VIN2 VDD GND VernierSymbol
x1 net3 net2 net4 net1 VDD GND VernierSymbol
x2 net5 net3 net6 net4 VDD GND VernierSymbol
x3 TEST1 net5 TEST2 net6 VDD GND VernierSymbol
x4 net8 TEST1 net7 TEST2 VDD GND VernierSymbol
x7 net9 net8 net10 net7 VDD GND VernierSymbol
x8 net11 net9 net12 net10 VDD GND VernierSymbol
x9 VOUT1 net11 VOUT2 net12 VDD GND VernierSymbol
**** begin user architecture code


.include $PDK_ROOT/sky130B/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.control
tran 10p 100n
write VernierDelay.raw
plot v(VOUT1) v(VOUT2) v(TEST1) V(TEST2)
.endc

.options acct list
.option numdgt=6


.lib /usr/local/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends

* expanding   symbol:  VernierSymbol.sym # of pins=6
** sym_path: /home/alexa/TemporalChip/xschem/projects/VernierSymbol.sym
** sch_path: /home/alexa/TemporalChip/xschem/projects/VernierSymbol.sch
.subckt VernierSymbol OUT1 IN1 OUT2 IN2 VDD GND
*.ipin VDD
*.ipin GND
*.ipin IN1
*.ipin IN2
*.opin OUT1
*.opin OUT2
x2 net8 OUT2 0 0 VDD VDD OUT1 sky130_fd_sc_hd__dlxtp_1
x10 net5 GND GND VDD VDD net7 sky130_fd_sc_hd__buf_1
x11 net4 GND GND VDD VDD net5 sky130_fd_sc_hd__buf_1
x12 IN2 GND GND VDD VDD net4 sky130_fd_sc_hd__buf_1
x6 net3 GND GND VDD VDD net6 sky130_fd_sc_hd__buf_1
x7 net2 GND GND VDD VDD net3 sky130_fd_sc_hd__buf_1
x8 net1 GND GND VDD VDD net2 sky130_fd_sc_hd__buf_1
x9 IN1 GND GND VDD VDD net1 sky130_fd_sc_hd__buf_1
x5 net6 GND GND VDD VDD net8 sky130_fd_sc_hd__buf_1
x13 net7 GND GND VDD VDD OUT2 sky130_fd_sc_hd__buf_1
.ends

.GLOBAL GND
.end
